* C:\Program Files\Orcad\Work\2015-2016-30-406\shemapokursovomubezkz.sch

* Schematics Version 9.2
* Wed Dec 02 07:30:29 2015



** Analysis setup **
.tran 0.1ms 25ms
.OPTIONS ABSTOL=100uA
.OPTIONS ITL4=40
.OPTIONS VNTOL=100uV
.LIB "C:\Program Files\Orcad\Work\2015-2016-30-406\Schematic1.lib"
.LIB "C:\Program Files\Orcad\Work\2015-2016-30-406\shemapokursovomubezkz.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "shemapokursovomubezkz.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
