* D:\GIT\MAI\viser\modeling\Start\SimmetrCM.sch

* Schematics Version 9.2
* Thu Mar 21 09:07:24 2019



** Analysis setup **
.tran 0ns 200m SKIPBP
.OPTIONS ABSTOL=1uA
.OPTIONS ITL4=70
.OPTIONS RELTOL=0.01


* From [PSPICE NETLIST] section of d:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "D:\Program Files\Orcad\PSpice\UserLib\OPA_2.lib"
.lib "D:\Program Files\Orcad\PSpice\UserLib\MyLib.lib"
.lib "nom.lib"

.INC "SimmetrCM.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
