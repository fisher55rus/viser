* D:\GIT\MAI\viser\modeling\220VDC\220vdc.sch

* Schematics Version 9.2
* Thu Mar 21 11:29:56 2019



** Analysis setup **
.tran 0ns 1 0 10u SKIPBP


* From [PSPICE NETLIST] section of d:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "D:\Program Files\Orcad\PSpice\UserLib\OPA_2.lib"
.lib "D:\Program Files\Orcad\PSpice\UserLib\MyLib.lib"
.lib "nom.lib"

.INC "220vdc.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
