* D:\GIT\MAI\viser\modeling\half_bridge\Shevcov\Nik\Sxema5IzmenitVuxod.sch

* Schematics Version 9.2
* Fri Mar 29 22:23:47 2019



** Analysis setup **
.tran 0 8ms 0 0.1ms
.OPTIONS ABSTOL=100u
.OPTIONS DIGINITSTATE=0
.OPTIONS ITL4=40
.OPTIONS VNTOL=100uV
.LIB "D:\GIT\MAI\viser\modeling\half_bridge\Shevcov\Vova_repalov_kurs_shev\Repalov\shemapokursovomubezkz.lib"


* From [PSPICE NETLIST] section of d:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "D:\Program Files\Orcad\PSpice\UserLib\OPA_2.lib"
.lib "D:\Program Files\Orcad\PSpice\UserLib\MyLib.lib"
.lib "nom.lib"

.INC "Sxema5IzmenitVuxod.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
